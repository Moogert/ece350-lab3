module lab3(in, out); 
	input in;
	output out; 
	assign out = in; 
	
endmodule 